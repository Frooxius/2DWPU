PLL40Mhz_inst : PLL40Mhz PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
