INT_SQRT_inst : INT_SQRT PORT MAP (
		radical	 => radical_sig,
		q	 => q_sig,
		remainder	 => remainder_sig
	);
